package org;
	
	type CPU {
		int cores;
		int threads;
		long clock;
		long cache;
		long fsb;
	}
	
	type FPGA {
		string family;
		string device;
		string package;
		string speed;
	}