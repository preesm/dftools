package epfl.stimm;

import org.stdio.ethernet.*;
import org.stdio.uart.*;
import org.units.*;
import org.memories.DDR2;
  
component compaq671b() {

	operator CPU T8300 {
		cores = 2;
		threads = 2 ;
		clock = 2.4 * 10^9;
		cache = 3 * 10**6;
		fsb = 800 * 10**6;
	}
	
	interface Ethernet eth0 {
		address = "192.168.1.10";
		port = 1024;
		type = EType.SOCK_STREAM;
	}
	
	interface Ethernet eth1 {
		address = "172.16.1.10";
		port = 1024;
	}
	
	interface Uart com1 {
		device = "COM1";
		//baudRate = EBaudrate.56700;
	}
	
	interface Uart com2 {
		device = "COM1";
		baudRate = 2;
	}
	
	memory DDR2 RAM {
		speed = 533 * 10**6;
		size = 4 * 10**9;
	}
	
}
