package epfl.stimm;

import org.stdio.*;
import org.units.*;
import org.memories.*;

device ml509() eth0, com1 {

	operator FPGA {
		family = "VIRTEX5";
		device = "xc5vlx110t";
		package = "ffg1136";
		speed = "1C";
	} V5;
	
	interface ethernet {
		address = "192.168.1.11";
		port = 1024;
	} <==> eth0;
	
	interface uart{
		device = "uart0";
		baudRate = EBaudrate.57600;
	} <==> com0;
	
	interface uart {
		device = "uart0";
		baudRate = EBaudrate.57600;
	} <==> com1;
	
	memory DDR2{
		speed = 400 * 10^6;
		size = 256 * 10^6;
	} ddr2pc4200;
	
	memory SRAM{
		speed := 200 * 10^6;
		size := 9 * 10^6;
	} ZBT;
	
};
	