package org.module;

library Memories {

	enum ERamType { DRAM, SRAM }
	
	class DDR2 {
		ERamType ramTyp = ERamType.DRAM;
		long size;
		long speed;
	}
	
	class SRAM {
		ERamType ramType = ERamType.SRAM;
		long size;
		long speed;
	}
	
}
	
	
	
