package org.stdio;

library uart {

	enum EBaudrate {
		110, 300, 600, 1200, 2400, 4800, 9600, 14400, 19200,
		38400, 56000, 57600, 115200, 128000, 256000 }

	// Data bits (5-8)
	enum EDataBits { 5, 6, 7, 8 }

	// Parity scheme
	enum EParity {
		NO_PARITY, ODD_PARITY, EVEN_PARITY,
		MARK_PARITY, SPACE_PARITY }

	// Stop bits
	enum EStopBits { ONE_STOP_BIT, ONE_5STOP_BITS, TWO_STOP_BITS }

	// Handshaking
	enum EHandshake { HandshakeOff, HandshakeHardware, HandshakeSoftware }

	// Definition of 
	class Uart {
		String device;
		EParity parity; //= NO_PARITY;
		EHandshake handShake;// = HandshakeOff;
		EStopBits stopBits;// = ONE_STOP_BIT;
		EDataBits dataBits;// = 8;
		EBaudrate baudRate;// = 9600;
	}

}