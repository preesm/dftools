package epfl.stimm;

import org.stdio.Ethernet.*;
import org.stdio.Uart.*;
import org.module.Units.*;
import org.module.Memories.*;

component Ml509 () {

	operator FPGA V5 {
		device = "xc5vlx110t";
		packaging = "ffg1136";
		speed = "1C";
	}
	
	interface Ethernet eth0_TEST {
		sockaddr.address = "192.168.1.11";
		sockaddr.port = 1024;
		sockaddr.addon.x = "Hello world!!!";
	}
	
	
	interface Uart com0 {
		device = "uart0";
		baudRate = EBaudrate.EBaud57600;
	}
	
	
	memory DDR2 ddr {
		speed = 10;
		size = 256 * 10;
	} 
	
	memory SRAM ZBT {
		speed = 200 * 10;
		size = 9 * (10 + 10);
	}
	
}