package epfl.stimm;

import org.stdio.ethernet.*;
import org.stdio.uart.*;
import org.units.*;
import org.memories.DDR2;
  
component compaq671b() /*eth0, eth1, com1, com2*/{

	operator CPU T8300 {
		// cores = 2;
		// threads = 2;
		// clock = 2.4 * 10^9;
		// cache = 3 * 10^6;
		// fsb = 800 * 10^6;
	}
	
	interface ethernet eth.eth0 <==> eth0 {
		// address = "192.168.1.10";
		// port = 1024;
	}
	
	interface ethernet eth.wifi <==> eth1 {
		// address = "172.16.1.10";
		// port = 1024;
	}
	
	interface uart com1 <==> com1 {
		// device = "COM1";
		// baudRate = EBaudrate.57600;
	}
	
	interface uart com4 <==> com2 {
		// device = "COM1";
		// baudRate = EB
	}
	
	memory DDR2 {
		// speed = 533 * 10^6;
		// size = 4 * 10^9;
	}
	
}
