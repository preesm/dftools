package epfl.stimm;

import org.stdio.*;
import org.units;
import org.memories.DDR2;
  
component compaq671b() /*eth0, eth1, com1, com2*/{

	T8300 : operator CPU {
		/*cores = 2;
		threads = 2;
		clock = 2.4 * 10^9;
		cache = 3 * 10^6;
		fsb = 800 * 10^6;*/
	} 
	
	eth.eth0 : interface ethernet <==> eth0 {
		/*address = "192.168.1.10";
		port = 1024;*/
	}
	
	eth.wifi : interface ethernet <==> eth1 {
		/*address = "172.16.1.10";
		port = 1024;*/
	}
	
	com1 : interface uart <==> com1 {
		/*device = "COM1";
		baudRate = EBaudrate.57600;*/
	}
	
	com4 : interface uart <==> com2 {
		/*device = "COM1";
		baudRate = EB*/
	}
	
	RAM : memory DDR2 {
		/*speed = 533 * 10^6;
		size = 4 * 10^9;*/
	}
	
}
