package org;

	enum ERamType { DRAM, SRAM };
	
	type {
		ERamType ramType = ERamType.DRAM;
		long size;
		long speed;
	} DDR2;
	
	type {
		ERamType ramType = ERamType.SDRAM;
		long size;
		long speed;
	} SRAM;