package org.module;

library Units {

	class CPU {
		int cores;
		int threads;  
		long clock;
		long cache;
		long fsb;
	}
	
	class FPGA {
		String family;
		String device;
		String packaging;
		String speed;
	}


}