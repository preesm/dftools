package org.stdio;

library Uart {

	enum EBaudrate {
		EBaud110, EBaud300, EBaud600, EBaud1200, EBaud2400, EBaud4800, EBaud9600,
		EBaud14400, EBaud19200, EBaud38400, EBaud56000, EBaud57600, EBaud115200, 
		EBaud128000, EBaud256000 }

	// Data bits (5-8)
	enum EDataBits { Data5, Data6, Data7, Data8 }

	// Parity scheme
	enum EParity {
		NO_PARITY, ODD_PARITY, EVEN_PARITY,
		MARK_PARITY, SPACE_PARITY }

	// Stop bits
	enum EStopBits { ONE_STOP_BIT, ONE_5STOP_BITS, TWO_STOP_BITS }

	// Handshaking
	enum EHandshake { HandshakeOff, HandshakeHardware, HandshakeSoftware }

	// Definition of 
	class Uart {
		String device;
		EParity parity = EParity.NO_PARITY;
		EHandshake handShake = EHandshake.HandshakeOff;
		EStopBits stopBits = EStopBits.ONE_STOP_BIT;
		EDataBits dataBits = EDataBits.Data8;
		EBaudrate baudRate = EBaudrate.EBaud9600;
	}

}